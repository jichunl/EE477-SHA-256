// This is the message scheduler module for SHA-256 accelerator which produces the Wt value for SHA-256 digest
//
module message scheduler
	(input 
	,input
	,output
	);

endmodule 
