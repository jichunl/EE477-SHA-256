// This is the pre-processing function for message scheduler and SHA-256_compression
// 
// input:
// 
// output:
//
module pre_processing (input [
