// This is the controller that communicates with FSB and multiple SHA256_cores
//
//
//
//
module SHA256_multicore
